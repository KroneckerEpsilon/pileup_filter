library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.STD_LOGIC_MATH.all;

package sipm is
	type sipmhit is 
		record
			v : integer;
		end record;
end package;
